module tb_processor();

    // add x3, x4, x2
    // 00000000001000100000000110110011

    logic clk;
    logic rst;

    processor dut
    (
        .clk ( clk ),
        .rst ( rst )
    );

    // clock generator
    initial
    begin
        clk = 0;
        forever
        begin
            #5 clk = 1;
            #5 clk = 0;
            // $display("pc: %b", dut.pc_out);

		    $display("pc_sel_br:%b", dut.br_taken);
		    $display("pc_sel_j:%b", dut.jump);

        end
    end

    // reset generator
    initial
    begin
        rst = 1;
        #10;
        rst = 0;
        #100;
        $display("Processor is running");
        $display("x1: %b", dut.reg_file_i.reg_mem[1]);
        $display("x2: %b", dut.reg_file_i.reg_mem[2]);
        $display("x1+x2-> x3: %b", dut.reg_file_i.reg_mem[3]);
        $display("loaded in x4: %b", dut.reg_file_i.reg_mem[4]);
        $display("loaded UI in x5: %b", dut.reg_file_i.reg_mem[5]);
        $display("loaded UI in x6: %b", dut.reg_file_i.reg_mem[6]);
        $finish;
    end

    // initialize memory
    initial
    begin
        $readmemh("inst.mem", dut.inst_mem_i.mem);
        $readmemb("rf.mem", dut.reg_file_i.reg_mem);
    end

    // dumping the waveform
    initial
    begin
        $dumpfile("processor.vcd");
        $dumpvars(0, dut);
    end

endmodule